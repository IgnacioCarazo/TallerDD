module maquina_cafe(input logic [3:0] btn, 
						  input logic [1:0] switch);


	reg[3:0] btn_seleccionado;


// falta el modulo sumador (N_BIT_ADDER)
// falta el modulo que guarda el monto total (REGISTER)

//sel_boton seleccionador_de_boton(btn, btn_seleccionado);

//ing_serving_time_module modulo_servido(btn_seleccionado, tiempo);

//drink_cost_module modulo_costo(btn_seleccionado, costo);

//falta el comparador de tiempos de servido (COUNTER Y COMPARATOR)

// falta el comparador de costo vs monto ingresado (COMPARATOR)


//FSM control(clk, rst, cancelar, btn, out); //cancelar es temporal




endmodule