
 //`timescale 1ns / 1ps  

module ALU_tb;

//Inputs
 reg[3:0] A,B;
 reg[3:0] ALU_Code;

//Outputs
 wire[3:0] ALU_Result;
 reg [3:0]flags;

 
 integer i;
 ALU test_unit(
				ALU_Code,
            A,B,                
            ALU_Result, 
            flags 
     );
    initial begin
	 
      A = 4'b0101;
      B = 4'b1001;
		
		/* 
		----------------------------------------------------------------------
		|ALU_Code|   ALU Operation
		----------------------------------------------------------------------
		| 0000  |   ALU_Out = A + B;
		----------------------------------------------------------------------
		| 0001  |   ALU_Out = A - B;
		----------------------------------------------------------------------
		| 0100  |   ALU_Out = A << 1;
		----------------------------------------------------------------------
		| 0101  |   ALU_Out = A >> 1;
		----------------------------------------------------------------------
		| 1000  |   ALU_Out = A and B;
		----------------------------------------------------------------------
		| 1001  |   ALU_Out = A or B;
		----------------------------------------------------------------------
		| 1010  |   ALU_Out = A xor B;
		----------------------------------------------------------------------*/
		
      ALU_Code = 4'b0000;
		#100;
		ALU_Code = 4'b0001;
		#100;
		ALU_Code = 4'b0100;
		#100;
		ALU_Code = 4'b0101;
		#100;
		ALU_Code = 4'b1000;
		#100;
		ALU_Code = 4'b1001;
		#100;
		ALU_Code = 4'b1010;
		#100;

      

      
    end
endmodule