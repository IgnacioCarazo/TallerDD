
 //`timescale 1ns / 1ps  

module ALU_tb;

//Inputs
 reg[3:0] A,B;
 reg[2:0] ALU_Code;

//Outputs
 reg[3:0] ALU_Result;
 
 //N,Z,C,V
 reg [3:0]flags;
 
 //display
 reg [6:0]display;
 
 
 ALU test_unit(
				ALU_Code,
            A,B,                
            ALU_Result, 
            flags,
				display
     );
    initial begin
	 		/* ALU Arithmetic and Logic Operations
		----------------------------------------------------------------------
		|ALU_Sel|   ALU Operation
		----------------------------------------------------------------------
		| 000  |   ALU_Out = A + B;
		----------------------------------------------------------------------
		| 001  |   ALU_Out = A - B;
		----------------------------------------------------------------------
		| 010  |   ALU_Out = A << 1;
		----------------------------------------------------------------------
		| 011  |   ALU_Out = A >> 1;
		----------------------------------------------------------------------
		| 100  |   ALU_Out = A and B;
		----------------------------------------------------------------------
		| 101  |   ALU_Out = A or B;
		----------------------------------------------------------------------
		| 110  |   ALU_Out = A xor B;
`		----------------------------------------------------------------------*/


	   flags = 4'b0000;
		
      A = 4'b0101;
      B = 4'b1001;
		
      ALU_Code = 3'b000;
		#100;
		ALU_Code = 3'b001;
		#100;
		ALU_Code = 3'b010;
		#100;
		ALU_Code = 3'b011;
		#100;
		ALU_Code = 3'b100;
		#100;
		ALU_Code = 3'b101;
		#100;
		ALU_Code = 3'b110;
		#100;
		
		A = 4'b1101;
      B = 4'b1101;
		
      ALU_Code = 3'b000;
		#100;
		ALU_Code = 3'b001;
		#100;
		ALU_Code = 3'b010;
		#100;
		ALU_Code = 3'b011;
		#100;
		ALU_Code = 3'b100;
		#100;
		ALU_Code = 3'b101;
		#100;
		ALU_Code = 3'b110;
		#100;
		
		A = 4'b1101;
      B = 4'b0001;
		
      ALU_Code = 3'b000;
		#100;
		ALU_Code = 3'b001;
		#100;
		ALU_Code = 3'b010;
		#100;
		ALU_Code = 3'b011;
		#100;
		ALU_Code = 3'b100;
		#100;
		ALU_Code = 3'b101;
		#100;
		ALU_Code = 3'b110;
		#100;
		
		A = 4'b0001;
      B = 4'b0000;
		
      ALU_Code = 3'b000;
		#100;
		ALU_Code = 3'b001;
		#100;
		ALU_Code = 3'b010;
		#100;
		ALU_Code = 3'b011;
		#100;
		ALU_Code = 3'b100;
		#100;
		ALU_Code = 3'b101;
		#100;
		ALU_Code = 3'b110;
		#100;

      

      
    end
endmodule