module ALU ();

	
	sumador hacersuma(A,B,tmp_adder,carry_adder);
	
endmodule