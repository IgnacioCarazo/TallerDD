module BitInput (input logic[0:7]bits)



endmodule